.SUBCKT CD4016B 1 2 3 4 5
* Specifications Harris data books
* 1 ANALOG INPUT
* 2 ANALOG OUTPUT
* 3 CONTROL
* 4 VDD (POSITIVE SUPPLY)
* 5 VSS (NEGATIVE SUPPLY)
*
RINP  3 11 1500
D1 11 4 D1
D2 5 11 D1
*
M1 12 11 4 4 MP4016A L=8U W=48U  AD=500P AS=500P PD=110U PS=110U
M2 12 11 5 5 MN4016A L=8U W=16U  AD=160P AS=160P PD=48U PS=48U
*
M1A 13 12 4 4 MP4016A L=8U W=96U  AD=500P AS=500P PD=110U PS=110U
M2A 13 12 5 5 MN4016A L=8U W=32U  AD=160P AS=160P PD=48U PS=48U
*
M3 1 12 2 4  MP4016A L=8U W=360U AD=3600P AS=3600P PD=900U PS=900U
M4 2 13 1 5  MN4016A L=8U W=120U AD=1080P AS=1080P PD=286U PS=286U
*
.MODEL MN4016A NMOS LEVEL=2 VTO=1.45 TOX=1000E-10 NSUB=4.7E16
+XJ=3U LD=2U UO=625 UCRIT=1E5 UEXP=0.45 UTRA=0.25 RD=15 RS=15 
+NEFF=2.5 VMAX=1E6 CGBO=3E-10 CGDO=10E-10 CGSO=10E-10 CJSW=2F
+NFS=4E12  GAMMA=2.2 LAMBDA=0.02
*
.MODEL MP4016A PMOS LEVEL=2 VTO=-1.5 TOX=1000E-10 NSUB=7.6E15
+XJ=3U LD=1.5U UO=225 UCRIT=3E5 UEXP=.5 UTRA=0.25 RD=15 RS=15
+NEFF=2.5 VMAX=1E5 CGBO=3E-10 CGDO=10E-10 CGSO=10E-10 CJSW=1F
+NFS=1E12  GAMMA=1.8 LAMBDA=0.02
* 
.MODEL D1 D IS=923.17E-18 RS=10 CJO=1.0000E-12 M=.3333  VJ=.75
+ ISR=100.00E-12  BV=35.357  IBV=10U  TT=5.0000E-9
.ENDS

